module kopt();
	reg a,b;
endmodule
