module minpool((logic clk,
          logic rst,
		  logic [7:0] ip_a, //input-
		  logic [7:0] ip_b, //logicb	
		  logic [7:0] ip_c, //logicc
		  logic [7:0] ip_d, //logicd
		  output reg signed [7:0] op, //output
          output reg PoolComplete);

endmodule